/***********************************************************
 *  Copyright (C) 2023 by JakodYuan (JakodYuan@outlook.com).
 *  All right reserved.
************************************************************/

package axi_env_pkg;
    import uvm_pkg::*;
    import svk_pkg::*;
    import svk_axi_pkg::*;

    `include "cust_axi_sys_env_cfg.sv"
    `include "axi_env.sv"


endpackage