/***********************************************************
 *  Copyright (C) 2023 by JakodYuan (JakodYuan@outlook.com).
 *  All right reserved.
************************************************************/

`include "tests/apb_base_test.sv"
`include "tests/apb_sanity.sv"
