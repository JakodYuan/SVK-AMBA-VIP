/***********************************************************
 *  Copyright (C) 2023 by JakodYuan (JakodYuan@outlook.com).
 *  All right reserved.
************************************************************/

`include "tests/axi_base_test.sv"
`include "tests/axi_sanity.sv"