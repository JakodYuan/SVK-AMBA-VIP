/***********************************************************
 *  Copyright (C) 2023 by JakodYuan (JakodYuan@outlook.com).
 *  All right reserved.
************************************************************/

`include "tests/ahb_base_test.sv"
`include "tests/ahb_sanity.sv"
