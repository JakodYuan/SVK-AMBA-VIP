/***********************************************************
 *  Copyright (C) 2023 by JakodYuan (JakodYuan@outlook.com).
 *  All right reserved.
************************************************************/

class cust_ahb_sys_env_cfg extends svk_ahb_sys_env_cfg;
    `uvm_object_utils(cust_ahb_sys_env_cfg)

    function new(string name="cust_ahb_sys_env_cfg");
        super.new(name);

        master_num = 1;
        slave_num  = 1;
        create_sub_cfg(master_num, slave_num);
        for(int i=0; i<master_num; ++i)begin
            master_cfg[i].work_mode                = svk_dec::MASTER;
            master_cfg[i].hready_time_out          = 1000;
            master_cfg[i].data_width               = 32;
            master_cfg[i].addr_width               = 32;
            master_cfg[i].enable_strb              = 1;
            master_cfg[i].cancle_after_error       = 1;
        end
        for(int i=0; i<slave_num; ++i)begin
            slave_cfg[i].work_mode                = svk_dec::SLAVE;
            slave_cfg[i].hready_time_out          = 1000;
            slave_cfg[i].data_width               = 32;
            slave_cfg[i].addr_width               = 32;
            slave_cfg[i].enable_strb              = 1;
            slave_cfg[i].cancle_after_error       = 1;
        end
    endfunction


endclass
