/***********************************************************
 *  Copyright (C) 2023 by JakodYuan (JakodYuan@outlook.com).
 *  All right reserved.
************************************************************/

package ahb_env_pkg;
    import uvm_pkg::*;
    import svk_pkg::*;
    import svk_ahb_pkg::*;

    `include "cust_ahb_sys_env_cfg.sv"
    `include "ahb_env.sv"


endpackage
