/***********************************************************
 *  Copyright (C) 2023 by JakodYuan (JakodYuan@outlook.com).
 *  All right reserved.
************************************************************/

package apb_env_pkg;
    import uvm_pkg::*;
    import svk_pkg::*;
    import svk_apb_pkg::*;

    `include "cust_apb_sys_env_cfg.sv"
    `include "apb_env.sv"


endpackage
